//Subject:     CO project 2 -Zero_Filled 
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      
//----------------------------------------------
//Date:        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Zero_Filled(
    data_i,
    data_o
    );
               
//I/O ports
input   [16-1:0] data_i;
output  [32-1:0] data_o;

//Internal Signals
reg     [32-1:0] data_o;
//Sign extended
always@(*)
begin
	data_o[31:16]<=data_i[15:0];
	data_o[15:0]<=0;
end
endmodule      
     
